/*
    CS/ECE 552 Spring '23
    Homework #2, Problem 2

    A multi-bit ALU module (defaults to 16-bit). It is designed to choose
    the correct operation to perform on 2 multi-bit numbers from rotate
    left, shift left, shift right arithmetic, shift right logical, add,
    or, xor, & and.  Upon doing this, it should output the multi-bit result
    of the operation, as well as drive the output signals Zero and Overflow
    (OFL).
*/
`default_nettype none
module alu (InA, InB, Cin, Oper, invA, invB, sign, Out, Zero, Ofl);

    parameter OPERAND_WIDTH = 16;    
    parameter NUM_OPERATIONS = 3;
       
    input wire  [OPERAND_WIDTH -1:0] InA ; // Input wire operand A
    input wire  [OPERAND_WIDTH -1:0] InB ; // Input wire operand B
    input wire                       Cin ; // Carry in
    input wire  [NUM_OPERATIONS-1:0] Oper; // Operation type
    input wire                       invA; // Signal to invert A
    input wire                       invB; // Signal to invert B
    input wire                       sign; // Signal for signed operation
    output wire [OPERAND_WIDTH -1:0] Out ; // Result of comput wireation
    output wire                      Ofl ; // Signal if overflow occured
    output wire                      Zero; // Signal if Out is 0

    /* YOUR CODE HERE */
//logic as follow:
//Opcode: 3'b000 shift_left A, ShAmt=B[3:0] 
//Opcode: 3'b001 shift_right_logical
//Opcode: 3'b010 rotate_left
//Opcode: 3'b011 shift_right_arith
//Opcode: 3'b100 A + B
//Opcode: 3'b101 A and B
//Opcode: 3'b110 A or B
//Opcode: 3'b111 A xor B

//inv A and inv B
wire [15:0] A,B;// the actually A, B which has been used in ALU
assign A=(invA)? ~InA : InA;
assign B=(invB)? ~InB : InB;

//result from shifter (000 to 011)
//module shifter (InBS, ShAmt, ShiftOper, OutBS);
wire [15:0] result_s;//result from shifter
shifter ALU_shifter(.OutBS(result_s), .InBS(A), .ShiftOper(Oper[1:0]), .ShAmt(B[3:0]));

//result from adder (100)
//module  cla16b(inA, inB, sum, cIn, cOut);
wire [15:0] result_a;//adder result
wire adder_cOut;// for unsign overflow test
cla16b ALU_adder(.sum(result_a), .cIn(Cin), .inA(A), .inB(B), .cOut(adder_cOut));

//result from and, or, xor (101,110,111)
wire [15:0] result_and, result_or, result_xor;
assign result_and = A & B;
assign result_or = A|B;
assign result_xor = A^B; 

//ALU logic
assign Out=(Oper[2]==1'b0)? result_s:
           (Oper==3'b100)? result_a:
           (Oper==3'b101)? result_and:
           (Oper==3'b110)? result_or:
           (Oper==3'b111)? result_xor : InA;

//Zero logic
assign Zero=(Out==16'd0)? 1'b1 : 1'b0;

//Overflow logic
//Only sign==1, there is an overflow
//
wire both_neg, both_pos;
wire Ofl_sign, Ofl_unsign;// for sign and unsign both need to test the over flow
assign both_neg=(A[15] & B[15])? 1'b1 : 1'b0;  
assign both_pos=((~A[15]) & (~B[15]))? 1'b1 : 1'b0; 
assign Ofl_sign=((both_neg) & (~Out[15])) | ((both_pos) & (Out[15]));
assign Ofl=(sign)? Ofl_sign: adder_cOut;

  
endmodule
`default_nettype wire
